`define RED       3'b100
`define GREEN     3'b010
`define BLUE      3'b001
`define BLACK     3'b000
`define WIGHT     3'b111
